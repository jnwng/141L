`timescale 1ns / 1ps

module pc
(
	input in,
	output reg out
);

always
begin
  out = in;
end

endmodule