library verilog;
use verilog.vl_types.all;
entity program_runner_2 is
end program_runner_2;
