library verilog;
use verilog.vl_types.all;
entity ALU_TB is
end ALU_TB;
