library verilog;
use verilog.vl_types.all;
entity NEXT_PC_TB is
end NEXT_PC_TB;
