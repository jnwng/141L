library verilog;
use verilog.vl_types.all;
entity program_runner_1 is
end program_runner_1;
