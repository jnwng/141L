library verilog;
use verilog.vl_types.all;
entity INSTR_ROM_TB is
end INSTR_ROM_TB;
